//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(148,144)(209,144){1}
//: {2}(213,144)(298,144){3}
//: {4}(211,146)(211,376)(366,376){5}
reg w1;    //: /sn:0 {0}(153,253)(180,253){1}
//: {2}(184,253)(283,253)(283,149)(298,149){3}
//: {4}(182,255)(182,381)(366,381){5}
reg w2;    //: /sn:0 {0}(149,333)(321,333)(321,319){1}
//: {2}(323,317)(375,317)(375,311)(390,311){3}
//: {4}(321,315)(321,152)(452,152){5}
wire w14;    //: /sn:0 {0}(473,150)(617,150)(617,138){1}
wire w3;    //: /sn:0 {0}(319,147)(366,147){1}
//: {2}(370,147)(452,147){3}
//: {4}(368,149)(368,306)(390,306){5}
wire w8;    //: /sn:0 {0}(387,379)(549,379)(549,314)(564,314){1}
wire w11;    //: /sn:0 {0}(585,312)(627,312)(627,300){1}
wire w5;    //: /sn:0 {0}(564,309)(411,309){1}
//: enddecls

  //: joint g8 (w0) @(211, 144) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g4 (.I0(w0), .I1(w1), .Z(w8));   //: @(377,379) /sn:0 /w:[ 5 5 0 ]
  //: LED g13 (w11) @(627,293) /sn:0 /w:[ 1 ] /type:0
  _GGAND2 #(6) g3 (.I0(w3), .I1(w2), .Z(w5));   //: @(401,309) /sn:0 /w:[ 5 3 1 ]
  //: SWITCH g2 (w2) @(132,333) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g1 (w1) @(136,253) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g11 (w2) @(321, 317) /w:[ 2 4 -1 1 ]
  //: joint g10 (w1) @(182, 253) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g6 (.I0(w3), .I1(w2), .Z(w14));   //: @(463,150) /sn:0 /w:[ 3 5 0 ]
  //: joint g9 (w3) @(368, 147) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g7 (.I0(w0), .I1(w1), .Z(w3));   //: @(309,147) /sn:0 /w:[ 3 3 0 ]
  _GGOR2 #(6) g5 (.I0(w5), .I1(w8), .Z(w11));   //: @(575,312) /sn:0 /w:[ 0 1 0 ]
  //: SWITCH g0 (w0) @(131,144) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: LED g12 (w14) @(617,131) /sn:0 /w:[ 1 ] /type:0

endmodule
//: /netlistEnd


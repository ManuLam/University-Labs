//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] w6;    //: /sn:0 {0}(696,213)(#:696,149){1}
supply0 w7;    //: /sn:0 {0}(436,138)(463,138)(463,164){1}
reg [7:0] w4;    //: /sn:0 {0}(571,211)(#:571,149){1}
reg w0;    //: /sn:0 {0}(73,155)(88,155){1}
reg [7:0] w31;    //: /sn:0 {0}(#:224,420)(224,405){1}
wire w32;    //: /sn:0 {0}(217,347)(217,362){1}
wire w16;    //: /sn:0 {0}(191,37)(206,37){1}
wire w14;    //: /sn:0 {0}(191,61)(206,61){1}
wire w19;    //: /sn:0 {0}(293,139)(293,124){1}
wire w15;    //: /sn:0 {0}(191,49)(206,49){1}
wire [7:0] w3;    //: /sn:0 {0}(412,219)(#:412,153){1}
wire [7:0] w34;    //: /sn:0 {0}(#:222,368)(222,383){1}
wire w21;    //: /sn:0 {0}(246,236)(246,221){1}
wire w28;    //: /sn:0 {0}(378,319)(393,319){1}
wire w24;    //: /sn:0 {0}(362,374)(362,359){1}
wire [1:0] w23;    //: /sn:0 {0}(#:320,337)(349,337){1}
wire w20;    //: /sn:0 {0}(283,139)(283,124){1}
wire [7:0] w1;    //: /sn:0 {0}(396,124)(396,78)(#:315,78)(315,162)(#:212,162){1}
wire w25;    //: /sn:0 {0}(378,355)(393,355){1}
wire [1:0] w18;    //: /sn:0 {0}(199,185)(199,200)(#:241,200)(#:241,215){1}
wire w8;    //: /sn:0 {0}(168,180)(183,180){1}
wire w30;    //: /sn:0 {0}(299,332)(314,332){1}
wire w22;    //: /sn:0 {0}(236,236)(236,221){1}
wire [1:0] w17;    //: /sn:0 {0}(222,78)(222,103)(#:288,103)(#:288,118){1}
wire w12;    //: /sn:0 {0}(168,144)(183,144){1}
wire w11;    //: /sn:0 {0}(168,156)(183,156){1}
wire [7:0] w2;    //: /sn:0 {0}(#:235,55)(428,55)(428,124){1}
wire w10;    //: /sn:0 {0}(168,168)(183,168){1}
wire w27;    //: /sn:0 {0}(378,331)(393,331){1}
wire w13;    //: /sn:0 {0}(191,73)(206,73){1}
wire w33;    //: /sn:0 {0}(227,347)(227,362){1}
wire w5;    //: /sn:0 {0}(339,110)(339,138)(388,138){1}
wire w29;    //: /sn:0 {0}(299,342)(314,342){1}
wire [7:0] w9;    //: /sn:0 {0}(#:412,235)(412,273){1}
//: {2}(414,275)(569,275){3}
//: {4}(573,275)(696,275)(#:696,229){5}
//: {6}(571,273)(#:571,227){7}
//: {8}(410,275)(342,275){9}
wire w26;    //: /sn:0 {0}(378,343)(393,343){1}
//: enddecls

  _GGBUF8 #(4) g8 (.I(w4), .Z(w9));   //: @(571,217) /sn:0 /R:3 /w:[ 0 7 ]
  //: DIP g4 (w4) @(571,139) /sn:0 /w:[ 1 ] /st:0 /dn:1
  tran g13[1:0] ({w19, w20}, w17);   //: @(288,119) /sn:0 /R:1 /dr:0 /tp:0 /drp:-1 /w:[ 1 1 1 ]
  //: GROUND g3 (w7) @(463,170) /sn:0 /w:[ 1 ]
  //: LED g2 (w5) @(339,103) /sn:0 /w:[ 0 ] /type:0
  _GGADD8 #(68, 70, 62, 64) g1 (.A(w1), .B(w2), .S(w3), .CI(w7), .CO(w5));   //: @(412,140) /sn:0 /w:[ 0 1 1 0 1 ]
  tran g16[1:0] ({w29, w30}, w23);   //: @(319,337) /sn:0 /dr:0 /tp:0 /drp:-1 /w:[ 1 1 0 ]
  _GGMUX4x8 #(12, 12) g11 (.I0(w8), .I1(w10), .I2(w11), .I3(w12), .S(w18), .Z(w1));   //: @(199,162) /sn:0 /R:1 /w:[ 1 1 1 1 0 1 ] /ss:0 /do:0
  //: joint g10 (w9) @(412, 275) /w:[ 2 1 8 -1 ]
  _GGBUF8 #(4) g6 (.I(w3), .Z(w9));   //: @(412,225) /sn:0 /R:3 /w:[ 0 0 ]
  //: joint g9 (w9) @(571, 275) /w:[ 4 6 3 -1 ]
  _GGBUF8 #(4) g7 (.I(w6), .Z(w9));   //: @(696,219) /sn:0 /R:3 /w:[ 0 5 ]
  _GGDECODER4 #(6, 6) g15 (.I(w23), .E(w24), .Z0(w25), .Z1(w26), .Z2(w27), .Z3(w28));   //: @(362,337) /sn:0 /R:1 /w:[ 1 1 0 0 0 0 ] /ss:0 /do:0
  //: DIP g17 (w31) @(224,431) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  tran g14[1:0] ({w21, w22}, w18);   //: @(241,216) /sn:0 /R:1 /dr:0 /tp:0 /drp:-1 /w:[ 1 1 1 ]
  //: DIP g5 (w6) @(696,139) /sn:0 /w:[ 1 ] /st:3 /dn:1
  //: SWITCH g0 (w0) @(56,155) /sn:0 /w:[ 0 ] /st:0 /dn:1
  tran g18[7:0] ({w32, w33}, w34);   //: @(222,367) /sn:0 /R:3 /dr:0 /tp:0 /drp:-1 /w:[ 1 1 0 ]
  _GGMUX4x8 #(12, 12) g12 (.I0(w13), .I1(w14), .I2(w15), .I3(w16), .S(w17), .Z(w2));   //: @(222,55) /sn:0 /R:1 /w:[ 1 1 1 1 0 0 ] /ss:0 /do:0

endmodule
//: /netlistEnd


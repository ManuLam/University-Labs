//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab10.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] w7;    //: /sn:0 {0}(#:647,677)(647,654)(647,654)(#:647,653){1}
reg w4;    //: /sn:0 {0}(301,81)(320,81)(320,171)(317,171){1}
//: {2}(313,171)(261,171){3}
//: {4}(315,173)(315,222)(341,222)(341,288){5}
//: {6}(339,290)(329,290)(329,293)(262,293){7}
//: {8}(341,292)(341,435){9}
//: {10}(339,437)(329,437)(329,438)(266,438){11}
//: {12}(341,439)(341,611)(255,611){13}
supply1 w19;    //: /sn:0 {0}(850,672)(850,623)(850,623)(850,608){1}
reg [7:0] w34;    //: /sn:0 {0}(1065,420)(#:1065,304){1}
supply0 w28;    //: /sn:0 {0}(881,310)(881,287)(860,287){1}
reg [7:0] w36;    //: /sn:0 {0}(1270,399)(1270,323)(#:1270,323)(#:1270,308){1}
reg w5;    //: /sn:0 {0}(509,720)(562,720)(562,231)(139,231)(139,216)(149,216){1}
//: {2}(153,216)(170,216)(170,176)(185,176){3}
//: {4}(151,218)(151,296){5}
//: {6}(153,298)(179,298)(179,298)(186,298){7}
//: {8}(151,300)(151,441){9}
//: {10}(153,443)(190,443){11}
//: {12}(151,445)(151,616)(179,616){13}
supply1 w9;    //: /sn:0 {0}(541,444)(541,445)(541,445)(541,430){1}
wire w32;    //: /sn:0 {0}(866,580)(1312,580)(1312,578){1}
//: {2}(1312,574)(1312,569){3}
//: {4}(1310,576)(1300,576)(1300,407)(1275,407){5}
wire [7:0] w6;    //: /sn:0 {0}(#:229,517)(238,517){1}
//: {2}(242,517)(284,517)(284,508){3}
//: {4}(240,515)(240,480)(241,480)(241,470){5}
//: {6}(243,468)(373,468)(373,189){7}
//: {8}(375,187)(453,187){9}
//: {10}(373,185)(373,57)(#:450,57){11}
//: {12}(239,468)(227,468)(#:227,454){13}
wire [7:0] w16;    //: /sn:0 {0}(#:453,175)(411,175)(411,173)(353,173){1}
//: {2}(351,171)(351,45)(450,45){3}
//: {4}(351,175)(351,725)(281,725){5}
//: {6}(279,723)(#:279,667){7}
//: {8}(277,725)(216,725)(#:216,627){9}
wire [7:0] w14;    //: /sn:0 {0}(852,273)(852,63)(#:479,63){1}
wire w15;    //: /sn:0 {0}(757,591)(612,591)(612,647){1}
wire [1:0] w3;    //: /sn:0 {0}(#:599,468)(569,468)(569,468)(554,468){1}
wire [7:0] w0;    //: /sn:0 {0}(#:267,365)(267,370)(223,370)(223,325){1}
//: {2}(225,323)(405,323)(405,200){3}
//: {4}(407,198)(#:417,198)(417,199)(453,199){5}
//: {6}(405,196)(405,69)(#:450,69){7}
//: {8}(223,321)(#:223,309){9}
wire w37;    //: /sn:0 {0}(758,264)(758,287)(812,287){1}
wire [7:0] w21;    //: /sn:0 {0}(#:482,193)(820,193)(820,273){1}
wire w31;    //: /sn:0 {0}(866,592)(1085,592)(1085,428)(1070,428){1}
wire [1:0] w20;    //: /sn:0 {0}(#:489,264)(469,264)(469,216){1}
wire w23;    //: /sn:0 {0}(495,269)(642,269)(642,647){1}
wire w24;    //: /sn:0 {0}(652,647)(652,387)(529,387)(529,134){1}
wire [7:0] w1;    //: /sn:0 {0}(#:1270,415)(1270,512)(1067,512){1}
//: {2}(1065,510)(#:1065,436){3}
//: {4}(1065,514)(1065,516)(838,516){5}
//: {6}(836,514)(#:836,389){7}
//: {8}(836,518)(836,528)(743,528)(743,568)(218,568){9}
//: {10}(214,568)(143,568)(143,420){11}
//: {12}(#:145,418)(227,418)(227,433){13}
//: {14}(143,416)(143,272){15}
//: {16}(#:145,270)(223,270)(223,288){17}
//: {18}(143,268)(143,133){19}
//: {20}(145,131)(222,131)(222,166){21}
//: {22}(141,131)(#:135,131){23}
//: {24}(216,570)(#:216,580)(216,580)(216,606){25}
wire w25;    //: /sn:0 {0}(539,134)(539,203)(662,203)(662,647){1}
wire w8;    //: /sn:0 {0}(525,462)(411,462)(411,303)(262,303){1}
wire w18;    //: /sn:0 {0}(255,621)(510,621)(510,486)(525,486){1}
wire [7:0] w35;    //: /sn:0 {0}(836,373)(836,319)(#:836,319)(#:836,302){1}
wire w30;    //: /sn:0 {0}(841,381)(912,381)(912,604)(866,604){1}
wire w17;    //: /sn:0 {0}(622,647)(622,581)(757,581){1}
wire w22;    //: /sn:0 {0}(495,259)(632,259)(632,647){1}
wire w2;    //: /sn:0 {0}(525,450)(440,450)(440,181)(261,181){1}
wire [1:0] w12;    //: /sn:0 {0}(466,86)(466,113)(#:534,113)(#:534,128){1}
wire [7:0] w10;    //: /sn:0 {0}(#:222,187)(222,216)(229,216){1}
//: {2}(233,216)(311,216)(311,197)(383,197){3}
//: {4}(387,197)(392,197)(392,211)(453,211){5}
//: {6}(385,195)(385,81)(450,81){7}
//: {8}(231,218)(231,236)(232,236)(232,242){9}
//: {10}(234,244)(277,244)(277,288)(307,288)(307,278){11}
//: {12}(230,244)(#:220,244){13}
wire w13;    //: /sn:0 {0}(266,448)(312,448)(312,474)(525,474){1}
wire w27;    //: /sn:0 {0}(605,473)(682,473)(682,647){1}
wire w33;    //: /sn:0 {0}(866,568)(881,568){1}
wire [1:0] w29;    //: /sn:0 {0}(837,586)(779,586)(#:779,586)(#:763,586){1}
wire w26;    //: /sn:0 {0}(605,463)(672,463)(672,647){1}
//: enddecls

  //: comment g4 @(220,258) /sn:0
  //: /line:"R1"
  //: /end
  //: comment g8 @(205,535) /sn:0
  //: /line:"R3"
  //: /end
  //: comment g3 @(222,103) /sn:0
  //: /line:"R0"
  //: /end
  //: joint g13 (w1) @(143, 131) /w:[ 20 -1 22 19 ]
  //: joint g34 (w0) @(405, 198) /w:[ 4 6 -1 3 ]
  _GGNDECODER4 #(4, 4) g37 (.I(w3), .E(w9), .Z0(w2), .Z1(w8), .Z2(w13), .Z3(w18));   //: @(541,468) /sn:0 /R:3 /w:[ 1 0 0 0 1 1 ] /ss:0 /do:0
  //: DIP g51 (w34) @(1065,294) /sn:0 /w:[ 1 ] /st:2 /dn:1
  _GGBUFIF8 #(4, 6) g55 (.Z(w1), .I(w36), .E(w32));   //: @(1270,405) /sn:0 /R:3 /w:[ 0 0 5 ]
  //: LED g58 (w10) @(307,271) /sn:0 /w:[ 11 ] /type:2
  _GGREG8 #(10, 10, 20) g2 (.Q(w0), .D(w1), .EN(w8), .CLR(w4), .CK(w5));   //: @(223,298) /sn:0 /w:[ 9 17 1 7 7 ]
  //: LED g59 (w0) @(267,358) /sn:0 /w:[ 0 ] /type:2
  //: SWITCH g1 (w5) @(492,720) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g16 (w1) @(216, 568) /w:[ 9 -1 10 24 ]
  //: joint g11 (w6) @(240, 517) /w:[ 2 4 1 -1 ]
  _GGBUFIF8 #(4, 6) g50 (.Z(w1), .I(w35), .E(w30));   //: @(836,379) /sn:0 /R:3 /w:[ 7 0 0 ]
  //: LED g10 (w6) @(284,501) /sn:0 /w:[ 3 ] /type:2
  //: joint g19 (w5) @(151, 443) /w:[ 10 9 -1 12 ]
  //: joint g32 (w6) @(373, 187) /w:[ 8 10 -1 7 ]
  _GGREG8 #(10, 10, 20) g6 (.Q(w16), .D(w1), .EN(w18), .CLR(w4), .CK(w5));   //: @(216,616) /sn:0 /w:[ 9 25 0 13 13 ]
  //: VDD g38 (w9) @(552,430) /sn:0 /w:[ 1 ]
  //: comment g7 @(224,368) /sn:0
  //: /line:"R2"
  //: /end
  //: joint g53 (w1) @(836, 516) /w:[ 5 6 -1 8 ]
  //: joint g57 (w32) @(1312, 576) /w:[ -1 2 4 1 ]
  //: joint g9 (w10) @(231, 216) /w:[ 2 -1 1 8 ]
  //: joint g15 (w1) @(143, 418) /w:[ 12 14 -1 11 ]
  //: comment g20 @(18,161) /sn:0
  //: /line:"Clock"
  //: /end
  //: joint g31 (w6) @(241, 468) /w:[ 6 -1 12 5 ]
  //: DIP g39 (w7) @(647,688) /sn:0 /R:2 /w:[ 0 ] /st:144 /dn:1
  assign w20 = {w23, w22}; //: CONCAT g43  @(490,264) /sn:0 /R:2 /w:[ 0 0 0 ] /dr:0 /tp:0 /drp:1
  //: LED g48 (w37) @(758,257) /sn:0 /w:[ 0 ] /type:0
  //: joint g17 (w5) @(151, 216) /w:[ 2 -1 1 4 ]
  //: joint g25 (w4) @(341, 437) /w:[ -1 9 10 12 ]
  _GGMUX4x8 #(12, 12) g29 (.I0(w10), .I1(w0), .I2(w6), .I3(w16), .S(w20), .Z(w21));   //: @(469,193) /sn:0 /R:1 /w:[ 5 5 9 0 1 0 ] /ss:0 /do:0
  assign w3 = {w27, w26}; //: CONCAT g42  @(600,468) /sn:0 /R:2 /w:[ 0 0 0 ] /dr:0 /tp:0 /drp:1
  _GGBUFIF8 #(4, 6) g52 (.Z(w1), .I(w34), .E(w31));   //: @(1065,426) /sn:0 /R:3 /w:[ 3 0 1 ]
  _GGREG8 #(10, 10, 20) g5 (.Q(w6), .D(w1), .EN(w13), .CLR(w4), .CK(w5));   //: @(227,443) /sn:0 /w:[ 13 13 0 11 11 ]
  //: joint g14 (w1) @(143, 270) /w:[ 16 18 -1 15 ]
  //: joint g56 (w1) @(1065, 512) /w:[ 1 2 -1 4 ]
  assign w29 = {w17, w15}; //: CONCAT g44  @(762,586) /sn:0 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:1
  _GGADD8 #(68, 70, 62, 64) g47 (.A(w21), .B(w14), .S(w35), .CI(w28), .CO(w37));   //: @(836,289) /sn:0 /w:[ 1 0 1 1 1 ]
  //: SWITCH g21 (w4) @(284,81) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: joint g24 (w4) @(341, 290) /w:[ -1 5 6 8 ]
  //: joint g36 (w10) @(385, 197) /w:[ 4 6 3 -1 ]
  //: joint g23 (w4) @(315, 171) /w:[ 1 -1 2 4 ]
  assign w12 = {w24, w25}; //: CONCAT g41  @(534,129) /sn:0 /R:1 /w:[ 1 1 0 ] /dr:0 /tp:0 /drp:1
  assign {w27, w26, w25, w24, w23, w22, w17, w15} = w7; //: CONCAT g40  @(647,652) /sn:0 /R:3 /w:[ 1 1 1 0 1 1 0 1 1 ] /dr:0 /tp:0 /drp:0
  //: DIP g54 (w36) @(1270,298) /sn:0 /w:[ 1 ] /st:2 /dn:1
  //: LED g60 (w16) @(279,660) /sn:0 /w:[ 7 ] /type:2
  _GGREG8 #(10, 10, 20) g0 (.Q(w10), .D(w1), .EN(w2), .CLR(w4), .CK(w5));   //: @(222,176) /sn:0 /w:[ 0 21 1 3 3 ]
  //: comment g22 @(269,22) /sn:0
  //: /line:"Clear"
  //: /line:"Registers"
  //: /end
  _GGMUX4x8 #(12, 12) g26 (.I0(w10), .I1(w0), .I2(w6), .I3(w16), .S(w12), .Z(w14));   //: @(466,63) /sn:0 /R:1 /w:[ 7 7 11 3 0 1 ] /ss:0 /do:0
  _GGDECODER4 #(6, 6) g45 (.I(w29), .E(w19), .Z0(w30), .Z1(w31), .Z2(w32), .Z3(w33));   //: @(850,586) /sn:0 /R:1 /w:[ 0 1 1 0 0 0 ] /ss:0 /do:0
  //: VDD g46 (w19) @(839,672) /sn:0 /R:2 /w:[ 0 ]
  //: joint g35 (w10) @(232, 244) /w:[ 10 9 12 -1 ]
  //: joint g18 (w5) @(151, 298) /w:[ 6 5 -1 8 ]
  //: joint g12 (w16) @(279, 725) /w:[ 5 6 8 -1 ]
  //: joint g30 (w16) @(351, 173) /w:[ 1 2 -1 4 ]
  //: joint g33 (w0) @(223, 323) /w:[ 2 8 -1 1 ]
  //: GROUND g49 (w28) @(881,316) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab5b.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(154,400)(196,400)(196,398){1}
//: {2}(198,396)(422,396)(422,252)(493,252){3}
//: {4}(196,394)(196,246)(211,246){5}
supply1 w12;    //: /sn:0 {0}(211,276)(87,276)(87,218){1}
//: {2}(89,216)(211,216){3}
//: {4}(87,214)(87,116){5}
reg w2;    //: /sn:0 {0}(306,327)(306,374){1}
//: {2}(308,376)(588,376)(588,333){3}
//: {4}(306,378)(306,444){5}
wire w4;    //: /sn:0 {0}(434,129)(434,156)(417,156)(417,226){1}
//: {2}(419,228)(443,228){3}
//: {4}(447,228)(478,228)(478,222)(493,222){5}
//: {6}(445,230)(445,282)(493,282){7}
//: {8}(415,228)(396,228){9}
wire [1:0] w1;    //: /sn:0 {0}(429,76)(#:429,123){1}
wire w11;    //: /sn:0 {0}(678,287)(693,287){1}
wire w10;    //: /sn:0 {0}(424,129)(424,151)(713,151)(713,234)(678,234){1}
wire w5;    //: /sn:0 {0}(396,281)(411,281){1}
//: enddecls

  //: SWITCH g4 (w0) @(137,400) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g8 (w4) @(417, 228) /w:[ 2 1 8 -1 ]
  //: joint g3 (w12) @(87, 216) /w:[ 2 4 -1 1 ]
  //: VDD g2 (w12) @(98,116) /sn:0 /w:[ 5 ]
  JKFlipFlop g1 (.K(w4), .CLK(w0), .J(w4), .RESET(w2), .Qinv(w11), .Q(w10));   //: @(494, 194) /sz:(183, 138) /sn:0 /p:[ Li0>7 Li1>3 Li2>5 Bi0>3 Ro0<0 Ro1<1 ]
  assign w1 = {w10, w4}; //: CONCAT g11  @(429,124) /sn:0 /R:1 /w:[ 1 0 0 ] /dr:0 /tp:0 /drp:1
  //: joint g10 (w4) @(445, 228) /w:[ 4 -1 3 6 ]
  //: joint g6 (w2) @(306, 376) /w:[ 2 1 -1 4 ]
  //: joint g9 (w0) @(196, 396) /w:[ 2 4 -1 1 ]
  //: LED g7 (w1) @(429,69) /sn:0 /w:[ 0 ] /type:3
  //: SWITCH g5 (w2) @(306,458) /sn:0 /R:1 /w:[ 5 ] /st:1 /dn:1
  JKFlipFlop g0 (.K(w12), .CLK(w0), .J(w12), .RESET(w2), .Qinv(w5), .Q(w4));   //: @(212, 188) /sz:(183, 138) /sn:0 /p:[ Li0>0 Li1>5 Li2>3 Bi0>0 Ro0<0 Ro1<9 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(CLK, K, Qinv, RESET, J, Q);
//: interface  /sz:(183, 138) /bd:[ Li0>K(88/138) Li1>CLK(58/138) Li2>J(28/138) Bi0>RESET(94/183) Ro0<Qinv(93/138) Ro1<Q(40/138) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(503,171)(520,171){1}
//: {2}(524,171)(573,171){3}
//: {4}(577,171)(671,171){5}
//: {6}(575,173)(575,252)(181,252)(181,210)(192,210){7}
//: {8}(522,173)(522,186)(541,186)(541,208)(470,208)(470,218)(480,218){9}
input K;    //: /sn:0 {0}(120,200)(192,200){1}
input J;    //: /sn:0 {0}(122,157)(197,157){1}
input RESET;    //: /sn:0 {0}(480,223)(271,223){1}
//: {2}(269,221)(269,215)(287,215){3}
//: {4}(269,225)(269,322){5}
output Qinv;    //: /sn:0 {0}(501,218)(521,218){1}
//: {2}(525,218)(546,218)(546,216)(593,216){3}
//: {4}(597,216)(669,216){5}
//: {6}(595,214)(595,118)(183,118)(183,167)(197,167){7}
//: {8}(523,216)(523,192)(468,192)(468,173)(482,173){9}
input CLK;    //: /sn:0 {0}(121,271)(154,271){1}
//: {2}(158,271)(195,271){3}
//: {4}(156,269)(156,207){5}
//: {6}(158,205)(192,205){7}
//: {8}(156,203)(156,162)(197,162){9}
//: {10}(156,273)(156,283)(171,283)(171,266)(195,266){11}
wire w20;    //: /sn:0 {0}(422,213)(480,213){1}
wire w8;    //: /sn:0 {0}(216,269)(367,269)(367,217){1}
//: {2}(369,215)(401,215){3}
//: {4}(367,213)(367,170)(400,170){5}
wire w17;    //: /sn:0 {0}(421,168)(482,168){1}
wire w2;    //: /sn:0 {0}(218,162)(285,162){1}
wire w11;    //: /sn:0 {0}(308,210)(323,210){1}
//: {2}(327,210)(401,210){3}
//: {4}(325,208)(325,183)(273,183)(273,167)(285,167){5}
wire w10;    //: /sn:0 {0}(306,165)(326,165){1}
//: {2}(330,165)(400,165){3}
//: {4}(328,167)(328,193)(276,193)(276,210)(287,210){5}
wire w5;    //: /sn:0 {0}(213,205)(287,205){1}
//: enddecls

  _GGNAND3 #(6) g4 (.I0(K), .I1(CLK), .I2(Q), .Z(w5));   //: @(203,205) /sn:0 /w:[ 1 7 7 0 ]
  _GGNAND2 #(4) g8 (.I0(w10), .I1(w8), .Z(w17));   //: @(411,168) /sn:0 /w:[ 3 5 0 ]
  _GGNAND3 #(6) g3 (.I0(J), .I1(CLK), .I2(Qinv), .Z(w2));   //: @(208,162) /sn:0 /w:[ 1 9 7 0 ]
  //: joint g13 (CLK) @(156, 205) /w:[ 6 8 -1 5 ]
  //: IN g2 (CLK) @(119,271) /sn:0 /w:[ 0 ]
  //: IN g1 (K) @(118,200) /sn:0 /w:[ 0 ]
  _GGNAND3 #(6) g11 (.I0(w20), .I1(Q), .I2(RESET), .Z(Qinv));   //: @(491,218) /sn:0 /w:[ 1 9 0 0 ]
  //: joint g16 (w8) @(367, 215) /w:[ 2 4 -1 1 ]
  _GGNAND2 #(4) g10 (.I0(w17), .I1(Qinv), .Z(Q));   //: @(493,171) /sn:0 /w:[ 1 9 0 ]
  //: OUT g19 (Qinv) @(666,216) /sn:0 /w:[ 5 ]
  _GGNAND3 #(6) g6 (.I0(w5), .I1(w10), .I2(RESET), .Z(w11));   //: @(298,210) /sn:0 /w:[ 1 5 3 0 ]
  _GGNAND2 #(4) g7 (.I0(w2), .I1(w11), .Z(w10));   //: @(296,165) /sn:0 /w:[ 1 5 0 ]
  _GGNAND2 #(4) g9 (.I0(w11), .I1(w8), .Z(w20));   //: @(412,213) /sn:0 /w:[ 3 3 0 ]
  //: joint g15 (w10) @(328, 165) /w:[ 2 -1 1 4 ]
  //: joint g20 (Qinv) @(595, 216) /w:[ 4 6 3 -1 ]
  //: joint g17 (w11) @(325, 210) /w:[ 2 4 1 -1 ]
  _GGNAND2 #(4) g5 (.I0(CLK), .I1(CLK), .Z(w8));   //: @(206,269) /sn:0 /w:[ 11 3 0 ]
  //: IN g14 (RESET) @(269,324) /sn:0 /R:1 /w:[ 5 ]
  //: joint g21 (Q) @(575, 171) /w:[ 4 -1 3 6 ]
  //: joint g24 (Qinv) @(523, 218) /w:[ 2 8 1 -1 ]
  //: joint g23 (Q) @(522, 171) /w:[ 2 -1 1 8 ]
  //: IN g0 (J) @(120,157) /sn:0 /w:[ 0 ]
  //: joint g22 (RESET) @(269, 223) /w:[ 1 2 -1 4 ]
  //: joint g12 (CLK) @(156, 271) /w:[ 2 4 1 10 ]
  //: OUT g18 (Q) @(668,171) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab5b.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(34,379)(134,379){1}
//: {2}(138,379)(420,379)(420,252)(493,252){3}
//: {4}(136,377)(136,242)(173,242){5}
reg w8;    //: /sn:0 {0}(106,269)(-12,269)(-12,216){1}
//: {2}(-10,214)(23,214){3}
//: {4}(27,214)(58,214){5}
//: {6}(25,212)(25,161)(365,161)(365,219)(395,219){7}
//: {8}(399,219)(446,219){9}
//: {10}(397,221)(397,282)(449,282){11}
//: {12}(-14,214)(-123,214){13}
reg w2;    //: /sn:0 {0}(268,458)(268,376)(268,376)(268,350){1}
//: {2}(270,348)(306,348)(306,364)(588,364)(588,333){3}
//: {4}(268,346)(268,323){5}
wire w6;    //: /sn:0 {0}(135,214)(74,214){1}
wire w7;    //: /sn:0 {0}(736,232)(759,232){1}
//: {2}(763,232)(784,232)(784,222){3}
//: {4}(761,230)(761,98)(103,98)(103,209)(135,209){5}
wire w16;    //: /sn:0 {0}(127,272)(173,272){1}
wire w4;    //: /sn:0 {0}(467,222)(493,222){1}
wire w1;    //: /sn:0 {0}(678,287)(736,287)(736,340)(82,340)(82,274)(106,274){1}
wire w18;    //: /sn:0 {0}(465,282)(493,282){1}
wire w12;    //: /sn:0 {0}(156,212)(173,212){1}
wire w10;    //: /sn:0 {0}(678,234)(715,234){1}
wire w5;    //: /sn:0 {0}(358,277)(373,277){1}
wire w9;    //: /sn:0 {0}(446,224)(424,224){1}
//: {2}(422,222)(422,155)(693,155)(693,229)(715,229){3}
//: {4}(420,224)(358,224){5}
//: enddecls

  //: comment g8 @(753,215) /sn:0
  //: /line:"Z"
  //: /end
  //: SWITCH g4 (w0) @(17,379) /sn:0 /w:[ 0 ] /st:1 /dn:1
  _GGOR2 #(6) g3 (.I0(w7), .I1(w6), .Z(w12));   //: @(146,212) /sn:0 /w:[ 5 0 0 ]
  _GGAND2 #(6) g13 (.I0(w8), .I1(w9), .Z(w4));   //: @(457,222) /sn:0 /w:[ 9 0 0 ]
  _GGNBUF #(2) g2 (.I(w8), .Z(w6));   //: @(64,214) /sn:0 /w:[ 5 1 ]
  JKFlipFlop g1 (.K(w18), .CLK(w0), .J(w4), .RESET(w2), .Qinv(w1), .Q(w10));   //: @(494, 194) /sz:(183, 138) /sn:0 /p:[ Li0>1 Li1>3 Li2>1 Bi0>3 Ro0<0 Ro1<0 ]
  //: joint g16 (w8) @(25, 214) /w:[ 4 6 3 -1 ]
  //: joint g11 (w9) @(422, 224) /w:[ 1 2 4 -1 ]
  //: joint g10 (w7) @(761, 232) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g19 (.I(w8), .Z(w18));   //: @(455,282) /sn:0 /w:[ 11 0 ]
  //: joint g6 (w2) @(268, 348) /w:[ 2 4 -1 1 ]
  //: comment g9 @(-78,186) /sn:0
  //: /line:"X"
  //: /end
  //: joint g7 (w0) @(136, 379) /w:[ 2 4 1 -1 ]
  //: LED g20 (w7) @(784,215) /sn:0 /w:[ 3 ] /type:0
  //: SWITCH g15 (w8) @(-140,214) /sn:0 /w:[ 13 ] /st:0 /dn:1
  //: joint g17 (w8) @(-12, 214) /w:[ 2 -1 12 1 ]
  _GGAND2 #(6) g14 (.I0(w8), .I1(w1), .Z(w16));   //: @(117,272) /sn:0 /w:[ 0 1 0 ]
  //: SWITCH g5 (w2) @(268,472) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  JKFlipFlop g0 (.K(w16), .CLK(w0), .J(w12), .RESET(w2), .Qinv(w5), .Q(w9));   //: @(174, 184) /sz:(183, 138) /sn:0 /p:[ Li0>1 Li1>5 Li2>1 Bi0>5 Ro0<0 Ro1<5 ]
  //: joint g18 (w8) @(397, 219) /w:[ 8 -1 7 10 ]
  _GGAND2 #(6) g12 (.I0(w9), .I1(w10), .Z(w7));   //: @(726,232) /sn:0 /w:[ 3 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin JKFlipFlop
module JKFlipFlop(CLK, K, Qinv, RESET, J, Q);
//: interface  /sz:(183, 138) /bd:[ Li0>J(28/138) Li1>CLK(58/138) Li2>K(88/138) Bi0>RESET(94/183) Ro0<Q(40/138) Ro1<Qinv(93/138) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(503,171)(520,171){1}
//: {2}(524,171)(573,171){3}
//: {4}(577,171)(671,171){5}
//: {6}(575,173)(575,252)(181,252)(181,210)(192,210){7}
//: {8}(522,173)(522,186)(541,186)(541,208)(470,208)(470,218)(480,218){9}
input K;    //: /sn:0 {0}(120,200)(192,200){1}
input RESET;    //: /sn:0 {0}(480,223)(271,223){1}
//: {2}(269,221)(269,215)(287,215){3}
//: {4}(269,225)(269,322){5}
input J;    //: /sn:0 {0}(122,157)(197,157){1}
output Qinv;    //: /sn:0 {0}(501,218)(521,218){1}
//: {2}(525,218)(546,218)(546,216)(593,216){3}
//: {4}(597,216)(669,216){5}
//: {6}(595,214)(595,118)(183,118)(183,167)(197,167){7}
//: {8}(523,216)(523,192)(468,192)(468,173)(482,173){9}
input CLK;    //: /sn:0 {0}(121,271)(154,271){1}
//: {2}(158,271)(195,271){3}
//: {4}(156,269)(156,207){5}
//: {6}(158,205)(192,205){7}
//: {8}(156,203)(156,162)(197,162){9}
//: {10}(156,273)(156,283)(171,283)(171,266)(195,266){11}
wire w20;    //: /sn:0 {0}(422,213)(480,213){1}
wire w8;    //: /sn:0 {0}(216,269)(367,269)(367,217){1}
//: {2}(369,215)(401,215){3}
//: {4}(367,213)(367,170)(400,170){5}
wire w17;    //: /sn:0 {0}(421,168)(482,168){1}
wire w11;    //: /sn:0 {0}(308,210)(323,210){1}
//: {2}(327,210)(401,210){3}
//: {4}(325,208)(325,183)(273,183)(273,167)(285,167){5}
wire w2;    //: /sn:0 {0}(218,162)(285,162){1}
wire w10;    //: /sn:0 {0}(306,165)(326,165){1}
//: {2}(330,165)(400,165){3}
//: {4}(328,167)(328,193)(276,193)(276,210)(287,210){5}
wire w5;    //: /sn:0 {0}(213,205)(287,205){1}
//: enddecls

  _GGNAND2 #(4) g8 (.I0(w10), .I1(w8), .Z(w17));   //: @(411,168) /sn:0 /w:[ 3 5 0 ]
  _GGNAND3 #(6) g4 (.I0(K), .I1(CLK), .I2(Q), .Z(w5));   //: @(203,205) /sn:0 /w:[ 1 7 7 0 ]
  //: joint g13 (CLK) @(156, 205) /w:[ 6 8 -1 5 ]
  _GGNAND3 #(6) g3 (.I0(J), .I1(CLK), .I2(Qinv), .Z(w2));   //: @(208,162) /sn:0 /w:[ 1 9 7 0 ]
  //: IN g2 (CLK) @(119,271) /sn:0 /w:[ 0 ]
  //: IN g1 (K) @(118,200) /sn:0 /w:[ 0 ]
  //: joint g16 (w8) @(367, 215) /w:[ 2 4 -1 1 ]
  _GGNAND3 #(6) g11 (.I0(w20), .I1(Q), .I2(RESET), .Z(Qinv));   //: @(491,218) /sn:0 /w:[ 1 9 0 0 ]
  _GGNAND2 #(4) g10 (.I0(w17), .I1(Qinv), .Z(Q));   //: @(493,171) /sn:0 /w:[ 1 9 0 ]
  //: OUT g19 (Qinv) @(666,216) /sn:0 /w:[ 5 ]
  _GGNAND3 #(6) g6 (.I0(w5), .I1(w10), .I2(RESET), .Z(w11));   //: @(298,210) /sn:0 /w:[ 1 5 3 0 ]
  _GGNAND2 #(4) g9 (.I0(w11), .I1(w8), .Z(w20));   //: @(412,213) /sn:0 /w:[ 3 3 0 ]
  _GGNAND2 #(4) g7 (.I0(w2), .I1(w11), .Z(w10));   //: @(296,165) /sn:0 /w:[ 1 5 0 ]
  //: joint g20 (Qinv) @(595, 216) /w:[ 4 6 3 -1 ]
  //: joint g15 (w10) @(328, 165) /w:[ 2 -1 1 4 ]
  //: joint g17 (w11) @(325, 210) /w:[ 2 4 1 -1 ]
  //: IN g14 (RESET) @(269,324) /sn:0 /R:1 /w:[ 5 ]
  _GGNAND2 #(4) g5 (.I0(CLK), .I1(CLK), .Z(w8));   //: @(206,269) /sn:0 /w:[ 11 3 0 ]
  //: joint g24 (Qinv) @(523, 218) /w:[ 2 8 1 -1 ]
  //: joint g21 (Q) @(575, 171) /w:[ 4 -1 3 6 ]
  //: joint g23 (Q) @(522, 171) /w:[ 2 -1 1 8 ]
  //: joint g22 (RESET) @(269, 223) /w:[ 1 2 -1 4 ]
  //: IN g0 (J) @(120,157) /sn:0 /w:[ 0 ]
  //: OUT g18 (Q) @(668,171) /sn:0 /w:[ 5 ]
  //: joint g12 (CLK) @(156, 271) /w:[ 2 4 1 10 ]

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab6.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 w3;    //: /sn:0 {0}(221,215)(185,215)(185,275)(192,275){1}
reg [3:0] w0;    //: /sn:0 {0}(#:80,305)(80,305)(80,305)(#:99,305){1}
reg [3:0] w1;    //: /sn:0 {0}(#:154,158)(154,156)(154,156)(#:154,202){1}
wire w6;    //: /sn:0 {0}(105,290)(139,290)(139,290)(192,290){1}
wire w7;    //: /sn:0 {0}(192,370)(129,370)(129,310)(105,310){1}
wire w14;    //: /sn:0 {0}(192,415)(124,415)(124,320)(105,320){1}
wire w15;    //: /sn:0 {0}(149,208)(149,383)(192,383){1}
wire w28;    //: /sn:0 {0}(192,339)(159,339)(159,208){1}
wire w23;    //: /sn:0 {0}(439,397)(529,397)(529,451){1}
wire w24;    //: /sn:0 {0}(439,358)(519,358)(519,451){1}
wire w25;    //: /sn:0 {0}(439,316)(509,316)(509,451){1}
wire w18;    //: /sn:0 {0}(105,300)(136,300)(136,328)(192,328){1}
wire w22;    //: /sn:0 {0}(439,425)(539,425)(539,451){1}
wire [4:0] w2;    //: /sn:0 {0}(#:519,457)(519,463)(616,463)(616,448){1}
wire w11;    //: /sn:0 {0}(192,426)(139,426)(139,208){1}
wire w27;    //: /sn:0 {0}(169,208)(169,261)(179,261)(179,301)(192,301){1}
wire w26;    //: /sn:0 {0}(439,283)(499,283)(499,451){1}
//: enddecls

  assign {w11, w15, w28, w27} = w1; //: CONCAT g4  @(154,203) /sn:0 /R:1 /w:[ 1 0 1 0 1 ] /dr:0 /tp:0 /drp:0
  assign {w14, w7, w18, w6} = w0; //: CONCAT g3  @(100,305) /sn:0 /R:2 /w:[ 1 1 0 0 1 ] /dr:0 /tp:0 /drp:0
  //: DIP g2 (w1) @(154,148) /sn:0 /w:[ 0 ] /st:0 /dn:1
  FourBitCarryLookAheadAdder g1 (.Cin(w3), .A0(w6), .B0(w27), .A1(w18), .B1(w28), .A2(w7), .B2(w15), .A3(w14), .B3(w11), .COUT0(w26), .COUT1(w25), .COUT2(w24), .COUT3(w23), .COUTall(w22));   //: @(193, 267) /sz:(245, 191) /sn:0 /p:[ Li0>1 Li1>1 Li2>1 Li3>1 Li4>0 Li5>0 Li6>1 Li7>0 Li8>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 ]
  assign w2 = {w22, w23, w24, w25, w26}; //: CONCAT g6  @(519,456) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  //: GROUND g7 (w3) @(227,215) /sn:0 /R:1 /w:[ 0 ]
  //: LED g5 (w2) @(616,441) /sn:0 /w:[ 1 ] /type:2
  //: DIP g0 (w0) @(42,305) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1

endmodule
//: /netlistEnd

//: /netlistBegin FourBitCarryLookAheadAdder
module FourBitCarryLookAheadAdder(A2, B1, A1, B0, A3, B3, B2, COUT0, COUT1, Cin, COUT3, COUT2, COUTall, A0);
//: interface  /sz:(245, 191) /bd:[ Li0>Cin(8/191) Li1>A0(23/191) Li2>B0(34/191) Li3>A1(61/191) Li4>B1(72/191) Li5>A2(103/191) Li6>B2(116/191) Li7>A3(148/191) Li8>B3(159/191) Ro0<COUT0(16/191) Ro1<COUT1(49/191) Ro2<COUT2(91/191) Ro3<COUT3(130/191) Ro4<COUTall(158/191) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input A0;    //: /sn:0 {0}(151,126)(141,126)(141,120)(127,120){1}
//: {2}(123,120)(117,120){3}
//: {4}(115,118)(115,100)(398,100){5}
//: {6}(113,120)(103,120){7}
//: {8}(125,122)(125,166)(152,166){9}
input A3;    //: /sn:0 {0}(127,422)(114,422)(114,413)(106,413){1}
//: {2}(102,413)(95,413){3}
//: {4}(91,413)(89,413){5}
//: {6}(93,415)(93,611)(391,611)(391,537)(457,537){7}
//: {8}(104,415)(104,455)(110,455){9}
//: {10}(114,455)(128,455){11}
//: {12}(112,457)(112,607)(385,607)(385,532)(457,532){13}
output COUTall;    //: /sn:0 {0}(457,542)(424,542)(424,515)(384,515){1}
//: {2}(382,513)(382,458)(504,458){3}
//: {4}(380,515)(349,515){5}
output COUT2;    //: /sn:0 {0}(419,210)(511,210){1}
input A2;    //: /sn:0 {0}(134,308)(121,308)(121,302)(111,302){1}
//: {2}(107,302)(100,302){3}
//: {4}(98,300)(98,290)(373,290)(373,324)(397,324){5}
//: {6}(96,302)(91,302){7}
//: {8}(109,304)(109,345)(136,345){9}
input B2;    //: /sn:0 {0}(92,322)(100,322){1}
//: {2}(104,322)(113,322){3}
//: {4}(117,322)(119,322)(119,313)(134,313){5}
//: {6}(115,320)(115,296)(365,296)(365,319)(397,319){7}
//: {8}(102,324)(102,350)(136,350){9}
input B1;    //: /sn:0 {0}(145,221)(128,221)(128,227)(125,227){1}
//: {2}(123,225)(123,205)(398,205){3}
//: {4}(121,227)(113,227){5}
//: {6}(109,227)(101,227){7}
//: {8}(111,229)(111,263)(145,263){9}
output COUT0;    //: /sn:0 {0}(419,105)(463,105)(463,105)(512,105){1}
output COUT1;    //: /sn:0 {0}(418,324)(506,324){1}
input Cin;    //: /sn:0 {0}(102,80)(219,80)(219,145){1}
//: {2}(221,147)(254,147){3}
//: {4}(219,149)(219,224){5}
//: {6}(221,226)(249,226){7}
//: {8}(219,228)(219,321){9}
//: {10}(221,323)(251,323){11}
//: {12}(219,325)(219,367)(219,367)(219,436){13}
//: {14}(221,438)(235,438)(235,438)(249,438){15}
//: {16}(219,440)(219,511){17}
input A1;    //: /sn:0 {0}(101,209)(107,209){1}
//: {2}(111,209)(115,209){3}
//: {4}(119,209)(132,209)(132,216)(145,216){5}
//: {6}(117,211)(117,258)(145,258){7}
//: {8}(109,207)(109,190)(373,190)(373,210)(398,210){9}
output COUT3;    //: /sn:0 {0}(478,537)(477,537)(477,537)(503,537){1}
input B3;    //: /sn:0 {0}(128,460)(98,460)(98,439){1}
//: {2}(100,437)(112,437)(112,427)(127,427){3}
//: {4}(96,437)(90,437){5}
input B0;    //: /sn:0 {0}(104,137)(107,137){1}
//: {2}(111,137)(114,137){3}
//: {4}(118,137)(141,137)(141,131)(151,131){5}
//: {6}(116,139)(116,171)(152,171){7}
//: {8}(109,135)(109,90)(366,90)(366,105)(398,105){9}
wire w6;    //: /sn:0 {0}(249,458)(171,458){1}
//: {2}(167,458)(149,458){3}
//: {4}(169,460)(169,501){5}
//: {6}(171,503)(247,503){7}
//: {8}(169,505)(169,552){9}
//: {10}(171,554)(247,554){11}
//: {12}(169,556)(169,586)(251,586){13}
wire w32;    //: /sn:0 {0}(344,359)(386,359)(386,329)(397,329){1}
wire w7;    //: /sn:0 {0}(275,150)(307,150){1}
wire w14;    //: /sn:0 {0}(328,510)(299,510)(299,448)(270,448){1}
wire w16;    //: /sn:0 {0}(269,276)(291,276)(291,247)(306,247){1}
wire w19;    //: /sn:0 {0}(323,357)(301,357)(301,330)(272,330){1}
wire w4;    //: /sn:0 {0}(247,544)(187,544)(187,398){1}
//: {2}(189,396)(251,396){3}
//: {4}(187,394)(187,221){5}
//: {6}(189,219)(191,219)(191,242)(306,242){7}
//: {8}(185,219)(166,219){9}
wire w0;    //: /sn:0 {0}(273,362)(323,362){1}
wire w3;    //: /sn:0 {0}(173,169)(206,169){1}
//: {2}(210,169)(239,169)(239,152)(254,152){3}
//: {4}(208,171)(208,229){5}
//: {6}(210,231)(249,231){7}
//: {8}(208,233)(208,326){9}
//: {10}(210,328)(251,328){11}
//: {12}(208,330)(208,441){13}
//: {14}(210,443)(249,443){15}
//: {16}(208,445)(208,521){17}
wire w31;    //: /sn:0 {0}(327,242)(386,242)(386,215)(398,215){1}
wire w1;    //: /sn:0 {0}(323,367)(274,367)(274,399)(272,399){1}
wire w25;    //: /sn:0 {0}(328,520)(277,520)(277,549)(268,549){1}
wire w18;    //: /sn:0 {0}(328,515)(277,515)(277,495)(268,495){1}
wire w8;    //: /sn:0 {0}(251,581)(175,581)(175,313){1}
//: {2}(177,311)(305,311)(305,352)(323,352){3}
//: {4}(173,311)(155,311){5}
wire w30;    //: /sn:0 {0}(328,148)(373,148)(373,110)(398,110){1}
wire w22;    //: /sn:0 {0}(272,584)(294,584)(294,525)(328,525){1}
wire w12;    //: /sn:0 {0}(270,231)(291,231)(291,237)(306,237){1}
wire w11;    //: /sn:0 {0}(148,425)(313,425)(313,505)(328,505){1}
wire w2;    //: /sn:0 {0}(172,129)(198,129){1}
//: {2}(202,129)(292,129)(292,145)(307,145){3}
//: {4}(200,131)(200,276){5}
//: {6}(202,278)(248,278){7}
//: {8}(200,280)(200,355){9}
//: {10}(202,357)(252,357){11}
//: {12}(200,359)(200,486){13}
//: {14}(202,488)(247,488){15}
//: {16}(200,490)(200,531){17}
wire w13;    //: /sn:0 {0}(166,261)(192,261){1}
//: {2}(196,261)(234,261)(234,236)(249,236){3}
//: {4}(194,263)(194,271){5}
//: {6}(196,273)(248,273){7}
//: {8}(194,275)(194,331){9}
//: {10}(196,333)(251,333){11}
//: {12}(194,335)(194,347)(194,347)(194,360){13}
//: {14}(196,362)(224,362)(224,362)(252,362){15}
//: {16}(194,364)(194,446){17}
//: {18}(196,448)(249,448){19}
//: {20}(194,450)(194,491){21}
//: {22}(196,493)(247,493){23}
//: {24}(194,495)(194,537){25}
wire w5;    //: /sn:0 {0}(247,549)(181,549)(181,500){1}
//: {2}(183,498)(247,498){3}
//: {4}(181,496)(181,455){5}
//: {6}(183,453)(249,453){7}
//: {8}(181,451)(181,403){9}
//: {10}(183,401)(251,401){11}
//: {12}(181,399)(181,369){13}
//: {14}(183,367)(252,367){15}
//: {16}(181,365)(181,340){17}
//: {18}(183,338)(251,338){19}
//: {20}(179,338)(172,338)(172,348)(157,348){21}
//: enddecls

  //: joint g61 (w4) @(187, 396) /w:[ 2 4 -1 1 ]
  _GGAND2 #(6) g8 (.I0(A0), .I1(B0), .Z(w2));   //: @(162,129) /sn:0 /w:[ 0 5 0 ]
  //: IN g4 (A2) @(89,302) /sn:0 /w:[ 7 ]
  //: joint g58 (w13) @(194, 362) /w:[ 14 13 -1 16 ]
  //: joint g55 (w3) @(208, 328) /w:[ 10 9 -1 12 ]
  //: joint g51 (w13) @(194, 273) /w:[ 6 5 -1 8 ]
  _GGOR2 #(6) g37 (.I0(w2), .I1(w7), .Z(w30));   //: @(318,148) /sn:0 /w:[ 3 1 0 ]
  _GGAND3 #(8) g34 (.I0(Cin), .I1(w3), .I2(w13), .Z(w12));   //: @(260,231) /sn:0 /w:[ 7 7 3 0 ]
  //: joint g13 (B0) @(116, 137) /w:[ 4 -1 3 6 ]
  //: IN g3 (B1) @(99,227) /sn:0 /w:[ 7 ]
  //: joint g86 (A3) @(112, 455) /w:[ 10 -1 9 12 ]
  //: joint g89 (B2) @(115, 322) /w:[ 4 6 3 -1 ]
  //: joint g77 (w6) @(169, 503) /w:[ 6 5 -1 8 ]
  //: joint g76 (w6) @(169, 458) /w:[ 1 -1 2 4 ]
  _GGAND4 #(10) g65 (.I0(w2), .I1(w13), .I2(w5), .I3(w6), .Z(w18));   //: @(258,495) /sn:0 /w:[ 15 23 3 7 1 ]
  //: IN g2 (A1) @(99,209) /sn:0 /w:[ 0 ]
  //: joint g59 (w5) @(181, 338) /w:[ 18 -1 20 17 ]
  //: joint g72 (w5) @(181, 453) /w:[ 6 8 -1 5 ]
  //: IN g1 (B0) @(102,137) /sn:0 /w:[ 0 ]
  _GGAND5 #(12) g64 (.I0(Cin), .I1(w3), .I2(w13), .I3(w5), .I4(w6), .Z(w14));   //: @(260,448) /sn:0 /w:[ 15 15 19 7 0 1 ]
  _GGXOR3 #(11) g98 (.I0(A0), .I1(B0), .I2(w30), .Z(COUT0));   //: @(409,105) /sn:0 /w:[ 5 9 1 0 ]
  _GGXOR3 #(11) g99 (.I0(A3), .I1(A3), .I2(COUTall), .Z(COUT3));   //: @(468,537) /sn:0 /w:[ 13 7 0 0 ]
  //: joint g16 (A1) @(117, 209) /w:[ 4 -1 3 6 ]
  _GGAND2 #(6) g11 (.I0(A3), .I1(B3), .Z(w11));   //: @(138,425) /sn:0 /w:[ 0 3 0 ]
  _GGXOR3 #(11) g96 (.I0(B2), .I1(A2), .I2(w32), .Z(COUT1));   //: @(408,324) /sn:0 /w:[ 7 5 1 0 ]
  //: joint g78 (w6) @(169, 554) /w:[ 10 9 -1 12 ]
  //: joint g50 (w4) @(187, 219) /w:[ 6 -1 8 5 ]
  //: comment g28 @(167,266) /sn:0
  //: /line:"P1"
  //: /end
  _GGAND2 #(6) g10 (.I0(A2), .I1(B2), .Z(w8));   //: @(145,311) /sn:0 /w:[ 0 5 5 ]
  //: joint g87 (A3) @(93, 413) /w:[ 3 -1 4 6 ]
  //: comment g32 @(153,467) /sn:0
  //: /line:"P3"
  //: /end
  //: comment g27 @(168,226) /sn:0
  //: /line:"G1"
  //: /end
  //: joint g19 (A2) @(109, 302) /w:[ 1 -1 2 8 ]
  //: joint g69 (w3) @(208, 443) /w:[ 14 13 -1 16 ]
  _GGOR3 #(8) g38 (.I0(w12), .I1(w4), .I2(w16), .Z(w31));   //: @(317,242) /sn:0 /w:[ 1 7 1 0 ]
  //: IN g6 (A3) @(87,413) /sn:0 /w:[ 5 ]
  //: joint g75 (w5) @(181, 498) /w:[ 2 4 -1 1 ]
  //: joint g57 (w2) @(200, 357) /w:[ 10 9 -1 12 ]
  _GGAND2 #(6) g53 (.I0(w4), .I1(w5), .Z(w1));   //: @(262,399) /sn:0 /w:[ 3 11 1 ]
  _GGOR2 #(6) g9 (.I0(A0), .I1(B0), .Z(w3));   //: @(163,169) /sn:0 /w:[ 9 7 0 ]
  //: IN g7 (B3) @(88,437) /sn:0 /w:[ 5 ]
  //: joint g71 (w8) @(175, 311) /w:[ 2 -1 4 1 ]
  //: comment g31 @(152,430) /sn:0
  //: /line:"G3"
  //: /end
  //: joint g20 (B2) @(102, 322) /w:[ 2 -1 1 8 ]
  _GGOR2 #(6) g15 (.I0(A1), .I1(B1), .Z(w13));   //: @(156,261) /sn:0 /w:[ 7 9 0 ]
  //: joint g68 (Cin) @(219, 438) /w:[ 14 13 -1 16 ]
  _GGAND3 #(8) g67 (.I0(w4), .I1(w5), .I2(w6), .Z(w25));   //: @(258,549) /sn:0 /w:[ 0 0 11 1 ]
  _GGOR4 #(10) g39 (.I0(w8), .I1(w19), .I2(w0), .I3(w1), .Z(w32));   //: @(334,359) /sn:0 /w:[ 3 0 1 0 0 ]
  //: joint g48 (w2) @(200, 278) /w:[ 6 5 -1 8 ]
  //: joint g43 (w3) @(208, 169) /w:[ 2 -1 1 4 ]
  //: joint g73 (w2) @(200, 488) /w:[ 14 13 -1 16 ]
  //: joint g62 (w5) @(181, 401) /w:[ 10 12 -1 9 ]
  //: comment g29 @(155,315) /sn:0
  //: /line:"G2"
  //: /end
  //: comment g25 @(173,135) /sn:0
  //: /line:"G0"
  //: /end
  //: joint g17 (B1) @(111, 227) /w:[ 5 -1 6 8 ]
  //: joint g88 (A2) @(98, 302) /w:[ 3 4 6 -1 ]
  _GGAND3 #(8) g52 (.I0(w2), .I1(w13), .I2(w5), .Z(w0));   //: @(263,362) /sn:0 /w:[ 11 15 15 0 ]
  //: comment g42 @(350,254) /sn:0
  //: /line:"Sum1"
  //: /end
  //: comment g63 @(361,530) /sn:0
  //: /line:"Sum3"
  //: /end
  //: joint g74 (w13) @(194, 493) /w:[ 22 21 -1 24 ]
  //: joint g56 (w13) @(194, 333) /w:[ 10 9 -1 12 ]
  _GGAND2 #(6) g14 (.I0(A1), .I1(B1), .Z(w4));   //: @(156,219) /sn:0 /w:[ 5 0 9 ]
  //: IN g5 (B2) @(90,322) /sn:0 /w:[ 0 ]
  _GGOR5 #(12) g79 (.I0(w11), .I1(w14), .I2(w18), .I3(w25), .I4(w22), .Z(COUTall));   //: @(339,515) /sn:0 /w:[ 1 0 0 0 1 5 ]
  //: joint g47 (w2) @(200, 129) /w:[ 2 -1 1 4 ]
  //: joint g44 (Cin) @(219, 226) /w:[ 6 5 -1 8 ]
  //: OUT g94 (COUT0) @(509,105) /sn:0 /w:[ 1 ]
  //: OUT g95 (COUT1) @(503,324) /sn:0 /w:[ 1 ]
  //: joint g80 (COUTall) @(382, 515) /w:[ 1 2 4 -1 ]
  _GGAND4 #(10) g36 (.I0(Cin), .I1(w3), .I2(w13), .I3(w5), .Z(w19));   //: @(262,330) /sn:0 /w:[ 11 11 11 19 1 ]
  //: IN g24 (Cin) @(100,80) /sn:0 /w:[ 0 ]
  _GGOR2 #(6) g21 (.I0(A3), .I1(B3), .Z(w6));   //: @(139,458) /sn:0 /w:[ 11 0 3 ]
  //: joint g84 (B0) @(109, 137) /w:[ 2 8 1 -1 ]
  //: joint g85 (A0) @(115, 120) /w:[ 3 4 6 -1 ]
  //: OUT g92 (COUT3) @(500,537) /sn:0 /w:[ 1 ]
  //: joint g23 (B3) @(98, 437) /w:[ 2 -1 4 1 ]
  //: comment g41 @(331,160) /sn:0
  //: /line:"Sum0"
  //: /end
  //: joint g60 (w5) @(181, 367) /w:[ 14 16 -1 13 ]
  //: joint g54 (Cin) @(219, 323) /w:[ 10 9 -1 12 ]
  //: joint g40 (Cin) @(219, 147) /w:[ 2 1 -1 4 ]
  //: OUT g93 (COUT2) @(508,210) /sn:0 /w:[ 1 ]
  //: OUT g81 (COUTall) @(501,458) /sn:0 /w:[ 3 ]
  //: joint g70 (w13) @(194, 448) /w:[ 18 17 -1 20 ]
  //: joint g45 (w3) @(208, 231) /w:[ 6 5 -1 8 ]
  _GGAND2 #(6) g35 (.I0(w13), .I1(w2), .Z(w16));   //: @(259,276) /sn:0 /w:[ 7 7 0 ]
  //: comment g26 @(174,175) /sn:0
  //: /line:"P0"
  //: /end
  //: joint g22 (A3) @(104, 413) /w:[ 1 -1 2 8 ]
  //: IN g0 (A0) @(101,120) /sn:0 /w:[ 7 ]
  //: comment g46 @(354,373) /sn:0
  //: /line:"Sum2"
  //: /end
  //: joint g90 (B1) @(123, 227) /w:[ 1 2 4 -1 ]
  _GGAND2 #(6) g66 (.I0(w8), .I1(w6), .Z(w22));   //: @(262,584) /sn:0 /w:[ 0 13 0 ]
  _GGXOR3 #(11) g97 (.I0(B1), .I1(A1), .I2(w31), .Z(COUT2));   //: @(409,210) /sn:0 /w:[ 3 9 1 0 ]
  _GGOR2 #(6) g18 (.I0(A2), .I1(B2), .Z(w5));   //: @(147,348) /sn:0 /w:[ 9 9 21 ]
  //: joint g12 (A0) @(125, 120) /w:[ 1 -1 2 8 ]
  _GGAND2 #(6) g33 (.I0(Cin), .I1(w3), .Z(w7));   //: @(265,150) /sn:0 /w:[ 3 3 0 ]
  //: comment g30 @(155,355) /sn:0
  //: /line:"P2"
  //: /end
  //: joint g91 (A1) @(109, 209) /w:[ 2 8 1 -1 ]
  //: joint g49 (w13) @(194, 261) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd


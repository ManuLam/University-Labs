//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab3B.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(-12,308)(-57,308)(-57,340)(-76,340){1}
reg w1;    //: /sn:0 {0}(406,166)(301,166)(301,245)(143,245){1}
reg a1;    //: /sn:0 {0}(314,374)(183,374)(183,256){1}
//: {2}(185,254)(316,254)(316,225)(378,225){3}
//: {4}(183,252)(183,186){5}
//: {6}(185,184)(264,184)(264,163)(278,163){7}
//: {8}(181,184)(94,184){9}
reg b1;    //: /sn:0 {0}(260,497)(200,497)(200,521)(172,521){1}
//: {2}(168,521)(157,521){3}
//: {4}(170,523)(170,620)(359,620){5}
reg a0;    //: /sn:0 {0}(314,369)(211,369)(211,146){1}
//: {2}(213,144)(264,144)(264,158)(278,158){3}
//: {4}(209,144)(142,144)(142,81)(110,81){5}
reg b0;    //: /sn:0 {0}(260,492)(199,492)(199,473)(187,473){1}
//: {2}(183,473)(155,473){3}
//: {4}(185,475)(185,615)(359,615){5}
reg w2;    //: /sn:0 {0}(-82,266)(-56,266)(-56,303)(-12,303){1}
wire w6;    //: /sn:0 {0}(19,374)(34,374){1}
wire w7;    //: /sn:0 {0}(50,374)(65,374){1}
wire w16;    //: /sn:0 {0}(453,573)(781,573)(781,377){1}
wire w14;    //: /sn:0 {0}(427,164)(703,164)(703,387)(718,387)(718,377){1}
wire w19;    //: /sn:0 {0}(363,257)(378,257){1}
wire w15;    //: /sn:0 {0}(380,618)(419,618)(419,575)(432,575){1}
wire w4;    //: /sn:0 {0}(391,500)(338,500){1}
//: {2}(334,500)(323,500)(323,447)(616,447)(616,312)(585,312){3}
//: {4}(336,502)(336,557)(354,557){5}
wire w3;    //: /sn:0 {0}(299,161)(367,161){1}
//: {2}(371,161)(406,161){3}
//: {4}(369,163)(369,220)(378,220){5}
wire w21;    //: /sn:0 {0}(340,576)(355,576){1}
wire w23;    //: /sn:0 {0}(376,579)(391,579){1}
wire w20;    //: /sn:0 {0}(399,255)(414,255){1}
wire w18;    //: /sn:0 {0}(363,252)(378,252){1}
wire w8;    //: /sn:0 {0}(335,372)(497,372)(497,314)(564,314){1}
wire w22;    //: /sn:0 {0}(340,581)(355,581){1}
wire w17;    //: /sn:0 {0}(48,409)(63,409){1}
wire w12;    //: /sn:0 {0}(412,498)(750,498)(750,377){1}
wire w11;    //: /sn:0 {0}(281,495)(308,495){1}
//: {2}(312,495)(391,495){3}
//: {4}(310,497)(310,552)(354,552){5}
wire w10;    //: /sn:0 {0}(17,409)(32,409){1}
wire w13;    //: /sn:0 {0}(375,555)(417,555)(417,570)(432,570){1}
wire w5;    //: /sn:0 {0}(564,309)(475,309)(475,223)(399,223){1}
wire w9;    //: /sn:0 {0}(9,306)(343,306){1}
//: {2}(345,304)(345,236){3}
//: {4}(345,308)(345,318)(290,318)(290,570){5}
//: enddecls

  //: joint g8 (a0) @(211, 144) /w:[ 2 -1 4 1 ]
  _GGAND2 #(6) g4 (.I0(a0), .I1(a1), .Z(w8));   //: @(325,372) /sn:0 /w:[ 0 0 0 ]
  _GGAND2 #(6) g37 (.I0(w18), .I1(w19), .Z(w20));   //: @(389,255) /sn:0 /w:[ 1 1 0 ]
  //: comment g34 @(773,342) /sn:0
  //: /line:"S2"
  //: /end
  //: SWITCH g13 (b0) @(138,473) /sn:0 /w:[ 3 ] /st:1 /dn:1
  _GGAND2 #(6) g3 (.I0(w3), .I1(a1), .Z(w5));   //: @(389,223) /sn:0 /w:[ 5 3 1 ]
  //: joint g2 (a1) @(183, 254) /w:[ 2 4 -1 1 ]
  //: SWITCH g1 (a1) @(77,184) /sn:0 /w:[ 9 ] /st:1 /dn:1
  //: SWITCH g11 (w2) @(-99,266) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGXOR2 #(8) g16 (.I0(w11), .I1(w4), .Z(w12));   //: @(402,498) /sn:0 /w:[ 3 0 0 ]
  //: SWITCH g28 (w0) @(-93,340) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: joint g10 (a1) @(183, 184) /w:[ 6 -1 8 5 ]
  //: comment g32 @(699,395) /sn:0
  //: /line:"Cout"
  //: /end
  //: joint g27 (w9) @(345, 306) /w:[ -1 2 1 4 ]
  //: joint g19 (w11) @(310, 495) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g38 (.I0(w21), .I1(w22), .Z(w23));   //: @(366,579) /sn:0 /w:[ 1 1 0 ]
  _GGXOR2 #(8) g6 (.I0(w3), .I1(w1), .Z(w14));   //: @(417,164) /sn:0 /w:[ 3 0 0 ]
  //: joint g9 (w3) @(369, 161) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g7 (.I0(a0), .I1(a1), .Z(w3));   //: @(289,161) /sn:0 /w:[ 3 7 0 ]
  //: comment g31 @(-152,340) /sn:0
  //: /line:"Sub"
  //: /end
  //: joint g20 (w4) @(336, 500) /w:[ 1 -1 2 4 ]
  _GGXOR2 #(8) g15 (.I0(b0), .I1(b1), .Z(w11));   //: @(271,495) /sn:0 /w:[ 0 0 0 ]
  //: SWITCH g29 (w1) @(126,245) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: LED g25 (w16) @(781,370) /sn:0 /w:[ 1 ] /type:0
  //: LED g17 (w12) @(750,370) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g14 (b1) @(140,521) /sn:0 /w:[ 3 ] /st:1 /dn:1
  _GGOR2 #(6) g5 (.I0(w5), .I1(w8), .Z(w4));   //: @(575,312) /sn:0 /w:[ 0 1 3 ]
  _GGNBUF #(2) g36 (.I(w10), .Z(w17));   //: @(38,409) /sn:0 /w:[ 1 0 ]
  _GGOR2 #(6) g24 (.I0(w13), .I1(w15), .Z(w16));   //: @(443,573) /sn:0 /w:[ 1 1 0 ]
  _GGAND2 #(6) g21 (.I0(b0), .I1(b1), .Z(w15));   //: @(370,618) /sn:0 /w:[ 5 5 0 ]
  //: joint g23 (b1) @(170, 521) /w:[ 1 -1 2 4 ]
  _GGNBUF #(2) g35 (.I(w6), .Z(w7));   //: @(40,374) /sn:0 /w:[ 1 0 ]
  _GGOR2 #(6) g26 (.I0(w2), .I1(w0), .Z(w9));   //: @(-1,306) /sn:0 /w:[ 1 0 0 ]
  //: joint g22 (b0) @(185, 473) /w:[ 1 -1 2 4 ]
  //: SWITCH g0 (a0) @(93,81) /sn:0 /w:[ 5 ] /st:1 /dn:1
  _GGAND2 #(6) g18 (.I0(w11), .I1(w4), .Z(w13));   //: @(365,555) /sn:0 /w:[ 5 5 0 ]
  //: LED g12 (w14) @(718,370) /sn:0 /w:[ 1 ] /type:0
  //: comment g33 @(744,342) /sn:0
  //: /line:"S1"
  //: /end
  //: comment g30 @(-153,259) /sn:0
  //: /line:"add"
  //: /end

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab4Aa.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w4;    //: /sn:0 {0}(177,464)(195,464){1}
//: {2}(199,464)(265,464){3}
//: {4}(197,466)(197,513)(215,513){5}
reg w0;    //: /sn:0 {0}(721,414)(690,414)(690,243)(702,243){1}
//: {2}(704,241)(704,165)(298,165){3}
//: {4}(296,163)(296,145)(233,145){5}
//: {6}(229,145)(219,145){7}
//: {8}(231,147)(231,277){9}
//: {10}(233,279)(274,279){11}
//: {12}(231,281)(231,415)(245,415)(245,518)(264,518){13}
//: {14}(296,167)(296,189)(332,189){15}
//: {16}(704,245)(704,348)(719,348){17}
reg w3;    //: /sn:0 {0}(182,364)(396,364){1}
reg w1;    //: /sn:0 {0}(332,194)(257,194){1}
//: {2}(253,194)(223,194){3}
//: {4}(255,196)(255,245){5}
//: {6}(257,247)(276,247){7}
//: {8}(255,249)(255,469)(265,469){9}
reg w2;    //: /sn:0 {0}(185,271)(197,271)(197,272){1}
//: {2}(199,274)(261,274)(261,252)(276,252){3}
//: {4}(197,276)(197,291)(212,291){5}
reg w5;    //: /sn:0 {0}(173,573)(382,573){1}
wire w6;    //: /sn:0 {0}(619,488)(550,488){1}
//: {2}(546,488)(481,488){3}
//: {4}(548,490)(548,533)(621,533){5}
wire w7;    //: /sn:0 {0}(228,291)(248,291)(248,284)(274,284){1}
wire w14;    //: /sn:0 {0}(640,491)(841,491){1}
wire w16;    //: /sn:0 {0}(740,351)(760,351)(760,336)(733,336)(733,295)(748,295){1}
wire w15;    //: /sn:0 {0}(295,282)(453,282)(453,266)(468,266){1}
wire w19;    //: /sn:0 {0}(669,358)(676,358){1}
//: {2}(680,358)(704,358)(704,353)(719,353){3}
//: {4}(678,360)(678,419)(721,419){5}
wire w34;    //: /sn:0 {0}(742,417)(1089,417)(1089,374){1}
wire w21;    //: /sn:0 {0}(769,293)(798,293)(798,511){1}
//: {2}(796,513)(784,513)(784,626)(803,626){3}
//: {4}(798,515)(798,543)(813,543){5}
wire w28;    //: /sn:0 {0}(841,496)(830,496)(830,510)(876,510)(876,546)(834,546){1}
wire w20;    //: /sn:0 {0}(417,367)(601,367){1}
//: {2}(605,367)(610,367)(610,292)(625,292){3}
//: {4}(603,365)(603,360)(648,360){5}
wire w24;    //: /sn:0 {0}(803,631)(753,631)(753,536)(751,536){1}
//: {2}(747,536)(642,536){3}
//: {4}(749,538)(749,548)(813,548){5}
wire w18;    //: /sn:0 {0}(619,493)(609,493)(609,494)(599,494){1}
//: {2}(595,494)(581,494)(581,571)(403,571){3}
//: {4}(597,496)(597,538)(621,538){5}
wire w8;    //: /sn:0 {0}(382,568)(372,568)(372,404){1}
//: {2}(374,402)(386,402)(386,369)(396,369){3}
//: {4}(372,400)(372,192)(353,192){5}
wire w35;    //: /sn:0 {0}(1157,443)(1157,629)(824,629){1}
wire w17;    //: /sn:0 {0}(285,516)(445,516)(445,490)(460,490){1}
wire w22;    //: /sn:0 {0}(646,290)(748,290){1}
wire w12;    //: /sn:0 {0}(286,467)(445,467)(445,485)(460,485){1}
wire w11;    //: /sn:0 {0}(297,250)(453,250)(453,261)(468,261){1}
wire w13;    //: /sn:0 {0}(489,264)(570,264){1}
//: {2}(574,264)(610,264)(610,287)(625,287){3}
//: {4}(572,266)(572,355)(648,355){5}
wire w29;    //: /sn:0 {0}(862,494)(1019,494)(1019,443){1}
wire w9;    //: /sn:0 {0}(231,513)(264,513){1}
//: enddecls

  //: SWITCH g4 (w4) @(160,464) /sn:0 /w:[ 0 ] /st:1 /dn:1
  _GGAND2 #(6) g8 (.I0(w4), .I1(w1), .Z(w12));   //: @(276,467) /sn:0 /w:[ 3 9 0 ]
  //: SWITCH g3 (w3) @(165,364) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g13 @(109,361) /sn:0
  //: /line:"A0"
  //: /end
  //: joint g34 (w18) @(597, 494) /w:[ 1 -1 2 4 ]
  //: joint g37 (w13) @(572, 264) /w:[ 2 -1 1 4 ]
  //: joint g51 (w0) @(704, 243) /w:[ -1 2 1 16 ]
  //: SWITCH g2 (w2) @(168,271) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g1 (w1) @(206,194) /sn:0 /w:[ 3 ] /st:0 /dn:1
  //: joint g11 (w4) @(197, 464) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g16 (.I0(w8), .I1(w5), .Z(w18));   //: @(393,571) /sn:0 /w:[ 0 1 3 ]
  _GGAND2 #(6) g10 (.I0(w9), .I1(w0), .Z(w17));   //: @(275,516) /sn:0 /w:[ 1 13 0 ]
  _GGAND2 #(6) g28 (.I0(w3), .I1(w8), .Z(w20));   //: @(407,367) /sn:0 /w:[ 1 3 0 ]
  //: joint g50 (w19) @(678, 358) /w:[ 2 -1 1 4 ]
  //: comment g19 @(162,185) /sn:0
  //: /line:"ADD"
  //: /end
  _GGOR2 #(6) g27 (.I0(w12), .I1(w17), .Z(w6));   //: @(471,488) /sn:0 /w:[ 1 1 3 ]
  _GGXOR2 #(8) g32 (.I0(w13), .I1(w20), .Z(w19));   //: @(659,358) /sn:0 /w:[ 5 5 0 ]
  _GGNBUF #(2) g6 (.I(w2), .Z(w7));   //: @(218,291) /sn:0 /w:[ 5 0 ]
  _GGOR2 #(6) g38 (.I0(w22), .I1(w16), .Z(w21));   //: @(759,293) /sn:0 /w:[ 1 1 0 ]
  _GGNBUF #(2) g7 (.I(w4), .Z(w9));   //: @(221,513) /sn:0 /w:[ 5 0 ]
  _GGAND2 #(6) g9 (.I0(w0), .I1(w7), .Z(w15));   //: @(285,282) /sn:0 /w:[ 11 1 0 ]
  //: comment g53 @(1093,342) /sn:0
  //: /line:"S1"
  //: /end
  //: comment g15 @(111,563) /sn:0
  //: /line:"A1"
  //: /end
  //: comment g20 @(162,138) /sn:0
  //: /line:"SUB"
  //: /end
  _GGAND2 #(6) g31 (.I0(w13), .I1(w20), .Z(w22));   //: @(636,290) /sn:0 /w:[ 3 3 0 ]
  _GGAND2 #(6) g39 (.I0(w0), .I1(w19), .Z(w16));   //: @(730,351) /sn:0 /w:[ 17 3 0 ]
  //: LED g43 (w34) @(1089,367) /sn:0 /w:[ 1 ] /type:0
  //: joint g48 (w0) @(296, 165) /w:[ 3 4 -1 14 ]
  _GGOR2 #(6) g17 (.I0(w0), .I1(w1), .Z(w8));   //: @(343,192) /sn:0 /w:[ 15 0 5 ]
  //: joint g25 (w1) @(255, 247) /w:[ 6 5 -1 8 ]
  //: joint g29 (w8) @(372, 402) /w:[ 2 4 -1 1 ]
  //: LED g42 (w29) @(1019,436) /sn:0 /w:[ 1 ] /type:0
  //: comment g52 @(1036,464) /sn:0
  //: /line:"Cout"
  //: /end
  //: SWITCH g5 (w5) @(156,573) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g14 @(109,456) /sn:0
  //: /line:"B1"
  //: /end
  //: LED g44 (w35) @(1157,436) /sn:0 /w:[ 0 ] /type:0
  //: joint g47 (w21) @(798, 513) /w:[ -1 1 2 4 ]
  //: joint g21 (w0) @(231, 145) /w:[ 5 -1 6 8 ]
  //: joint g24 (w2) @(197, 274) /w:[ 2 1 -1 4 ]
  //: joint g36 (w20) @(603, 367) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g23 (.I0(w1), .I1(w2), .Z(w11));   //: @(287,250) /sn:0 /w:[ 7 3 0 ]
  _GGAND2 #(6) g41 (.I0(w21), .I1(w24), .Z(w28));   //: @(824,546) /sn:0 /w:[ 5 5 1 ]
  _GGOR2 #(6) g40 (.I0(w14), .I1(w28), .Z(w29));   //: @(852,494) /sn:0 /w:[ 1 0 0 ]
  //: comment g54 @(1189,438) /sn:0
  //: /line:"S0"
  //: /end
  //: SWITCH g0 (w0) @(202,145) /sn:0 /w:[ 7 ] /st:1 /dn:1
  //: joint g22 (w0) @(231, 279) /w:[ 10 9 -1 12 ]
  _GGOR2 #(6) g26 (.I0(w11), .I1(w15), .Z(w13));   //: @(479,264) /sn:0 /w:[ 1 1 0 ]
  //: joint g35 (w6) @(548, 488) /w:[ 1 -1 2 4 ]
  _GGXOR2 #(8) g45 (.I0(w21), .I1(w24), .Z(w35));   //: @(814,629) /sn:0 /w:[ 3 0 1 ]
  //: joint g46 (w24) @(749, 536) /w:[ 1 -1 2 4 ]
  //: comment g12 @(108,252) /sn:0
  //: /line:"B0"
  //: /end
  //: joint g18 (w1) @(255, 194) /w:[ 1 -1 2 4 ]
  _GGAND2 #(6) g30 (.I0(w6), .I1(w18), .Z(w14));   //: @(630,491) /sn:0 /w:[ 0 0 0 ]
  _GGXOR2 #(8) g33 (.I0(w6), .I1(w18), .Z(w24));   //: @(632,536) /sn:0 /w:[ 5 5 3 ]
  _GGXOR2 #(8) g49 (.I0(w0), .I1(w19), .Z(w34));   //: @(732,417) /sn:0 /w:[ 0 5 0 ]

endmodule
//: /netlistEnd


//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply1 w6;    //: /sn:0 {0}(345,170)(316,170)(316,182){1}
//: {2}(318,184)(345,184){3}
//: {4}(316,186)(316,261){5}
supply0 w4;    //: /sn:0 {0}(345,150)(260,150)(260,175){1}
//: {2}(262,177)(345,177){3}
//: {4}(260,179)(260,185)(261,185)(261,188){5}
//: {6}(263,190)(345,190){7}
//: {8}(261,192)(261,261){9}
reg w3;    //: /sn:0 {0}(361,356)(361,264){1}
reg w0;    //: /sn:0 {0}(161,197)(218,197){1}
reg w1;    //: /sn:0 {0}(351,264)(351,340)(288,340)(288,355){1}
reg w2;    //: /sn:0 {0}(371,264)(371,341)(424,341)(424,356){1}
wire w16;    //: /sn:0 {0}(374,174)(430,174){1}
wire [2:0] w15;    //: /sn:0 {0}(#:361,258)(361,197){1}
wire w5;    //: /sn:0 {0}(234,197)(292,197){1}
//: {2}(296,197)(345,197){3}
//: {4}(294,195)(294,166){5}
//: {6}(296,164)(345,164){7}
//: {8}(294,162)(294,157)(345,157){9}
//: enddecls

  //: joint g8 (w5) @(294, 197) /w:[ 2 4 1 -1 ]
  _GGNBUF #(2) g4 (.I(w0), .Z(w5));   //: @(224,197) /sn:0 /w:[ 1 0 ]
  //: joint g13 (w6) @(316, 184) /w:[ 2 1 -1 4 ]
  //: SWITCH g3 (w3) @(361,370) /sn:0 /R:1 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g2 (w2) @(424,370) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g1 (w1) @(288,369) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  //: comment g16 @(360,394) /sn:0 /R:2
  //: /line:"B"
  //: /end
  //: LED g11 (w16) @(437,174) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g10 (w4) @(261, 190) /w:[ 6 5 -1 8 ]
  //: VDD g6 (w6) @(305,261) /sn:0 /R:2 /w:[ 5 ]
  //: joint g9 (w5) @(294, 164) /w:[ 6 8 -1 5 ]
  _GGMUX8 #(20, 20) g7 (.I0(w5), .I1(w4), .I2(w6), .I3(w4), .I4(w6), .I5(w5), .I6(w5), .I7(w4), .S(w15), .Z(w16));   //: @(361,174) /sn:0 /R:1 /w:[ 3 7 3 3 0 7 9 0 1 0 ] /ss:0 /do:0
  //: comment g15 @(418,396) /sn:0 /R:2
  //: /line:"A"
  //: /end
  //: comment g17 @(287,392) /sn:0 /R:2
  //: /line:"C"
  //: /end
  assign w15 = {w2, w3, w1}; //: CONCAT g14  @(361,259) /sn:0 /R:1 /w:[ 0 0 1 0 ] /dr:1 /tp:0 /drp:1
  //: GROUND g5 (w4) @(261,267) /sn:0 /w:[ 9 ]
  //: SWITCH g0 (w0) @(144,197) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g12 (w4) @(260, 177) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd


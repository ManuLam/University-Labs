//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Lab2LT.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(110,132)(195,132){1}
reg w3;    //: /sn:0 {0}(282,340)(231,340){1}
//: {2}(229,338)(229,236)(280,236){3}
//: {4}(229,342)(229,430)(110,430){5}
reg w1;    //: /sn:0 {0}(192,231)(109,231){1}
reg w2;    //: /sn:0 {0}(271,167)(153,167)(153,341)(129,341){1}
//: {2}(127,339)(127,335)(282,335){3}
//: {4}(125,341)(107,341){5}
wire w7;    //: /sn:0 {0}(208,231)(222,231){1}
//: {2}(226,231)(280,231){3}
//: {4}(224,233)(224,330)(282,330){5}
wire w16;    //: /sn:0 {0}(382,248)(319,248)(319,231)(301,231){1}
wire w19;    //: /sn:0 {0}(382,253)(331,253)(331,335)(303,335){1}
wire w8;    //: /sn:0 {0}(403,248)(468,248)(468,237){1}
wire w13;    //: /sn:0 {0}(382,243)(340,243)(340,165)(292,165){1}
wire w5;    //: /sn:0 {0}(280,226)(231,226)(231,134){1}
//: {2}(233,132)(256,132)(256,162)(271,162){3}
//: {4}(229,132)(211,132){5}
//: enddecls

  _GGNBUF #(2) g4 (.I(w0), .Z(w5));   //: @(201,132) /sn:0 /w:[ 1 5 ]
  _GGAND3 #(8) g8 (.I0(w5), .I1(w7), .I2(w3), .Z(w16));   //: @(291,231) /sn:0 /w:[ 0 3 3 1 ]
  //: SWITCH g3 (w3) @(93,430) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: joint g13 (w3) @(229, 340) /w:[ 1 2 -1 4 ]
  //: SWITCH g2 (w2) @(90,341) /sn:0 /w:[ 5 ] /st:1 /dn:1
  //: SWITCH g1 (w1) @(92,231) /sn:0 /w:[ 1 ] /st:1 /dn:1
  //: joint g11 (w7) @(224, 231) /w:[ 2 -1 1 4 ]
  //: joint g10 (w5) @(231, 132) /w:[ 2 -1 4 1 ]
  _GGOR3 #(8) g6 (.I0(w13), .I1(w16), .I2(w19), .Z(w8));   //: @(393,248) /sn:0 /w:[ 0 0 0 0 ]
  _GGAND2 #(6) g7 (.I0(w5), .I1(w2), .Z(w13));   //: @(282,165) /sn:0 /w:[ 3 0 1 ]
  _GGAND3 #(8) g9 (.I0(w7), .I1(w2), .I2(w3), .Z(w19));   //: @(293,335) /sn:0 /w:[ 5 3 0 1 ]
  _GGNBUF #(2) g5 (.I(w1), .Z(w7));   //: @(198,231) /sn:0 /w:[ 0 0 ]
  //: LED g14 (w8) @(468,230) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g0 (w0) @(93,132) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g12 (w2) @(127, 341) /w:[ 1 2 4 -1 ]

endmodule
//: /netlistEnd


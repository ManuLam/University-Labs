//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w3;    //: /sn:0 {0}(105,348)(160,348){1}
reg w0;    //: /sn:0 {0}(312,334)(268,334)(268,108)(161,108){1}
//: {2}(157,108)(100,108){3}
//: {4}(159,110)(159,114)(312,114){5}
reg w1;    //: /sn:0 {0}(104,186)(120,186){1}
//: {2}(122,184)(122,177)(315,177){3}
//: {4}(122,188)(122,339)(312,339){5}
reg w2;    //: /sn:0 {0}(105,272)(166,272){1}
wire w7;    //: /sn:0 {0}(315,182)(227,182)(227,346){1}
//: {2}(229,348)(299,348)(299,344)(312,344){3}
//: {4}(225,348)(176,348){5}
wire w15;    //: /sn:0 {0}(333,339)(420,339)(420,229)(435,229){1}
wire w4;    //: /sn:0 {0}(456,229)(563,229)(563,216){1}
wire w12;    //: /sn:0 {0}(435,234)(351,234)(351,177)(336,177){1}
wire w5;    //: /sn:0 {0}(315,172)(214,172)(214,272)(199,272){1}
//: {2}(197,270)(197,119)(312,119){3}
//: {4}(195,272)(182,272){5}
wire w9;    //: /sn:0 {0}(435,224)(406,224)(406,117)(333,117){1}
//: enddecls

  _GGAND3 #(8) g8 (.I0(w5), .I1(w1), .I2(w7), .Z(w12));   //: @(326,177) /sn:0 /w:[ 0 3 0 1 ]
  _GGNBUF #(2) g4 (.I(w2), .Z(w5));   //: @(172,272) /sn:0 /w:[ 1 5 ]
  //: joint g13 (w0) @(159, 108) /w:[ 1 -1 2 4 ]
  //: SWITCH g3 (w3) @(88,348) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g2 (w2) @(88,272) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g1 (w1) @(87,186) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g11 (w7) @(227, 348) /w:[ 2 1 4 -1 ]
  //: joint g10 (w1) @(122, 186) /w:[ -1 2 1 4 ]
  _GGNBUF #(2) g6 (.I(w3), .Z(w7));   //: @(166,348) /sn:0 /w:[ 1 5 ]
  _GGAND3 #(8) g9 (.I0(w0), .I1(w1), .I2(w7), .Z(w15));   //: @(323,339) /sn:0 /w:[ 0 5 3 0 ]
  _GGAND2 #(6) g7 (.I0(w0), .I1(w5), .Z(w9));   //: @(323,117) /sn:0 /w:[ 5 3 1 ]
  _GGOR3 #(8) g14 (.I0(w9), .I1(w15), .I2(w12), .Z(w4));   //: @(446,229) /sn:0 /w:[ 0 1 0 0 ]
  //: LED g5 (w4) @(563,209) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g0 (w0) @(83,108) /sn:0 /w:[ 3 ] /st:0 /dn:1
  //: joint g12 (w5) @(197, 272) /w:[ 1 2 4 -1 ]

endmodule
//: /netlistEnd


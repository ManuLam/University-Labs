//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "new.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg b;    //: /sn:0 {0}(47,207)(89,207){1}
//: {2}(93,207)(144,207){3}
//: {4}(91,205)(91,180){5}
//: {6}(93,178)(231,178)(231,177)(368,177){7}
//: {8}(91,176)(91,39)(363,39){9}
reg d;    //: /sn:0 {0}(368,187)(74,187){1}
//: {2}(72,185)(72,49)(363,49){3}
//: {4}(72,189)(72,354){5}
//: {6}(74,356)(141,356){7}
//: {8}(70,356)(49,356){9}
reg a;    //: /sn:0 {0}(367,277)(286,277)(286,261)(100,261)(100,141){1}
//: {2}(102,139)(110,139){3}
//: {4}(114,139)(142,139){5}
//: {6}(112,137)(112,34)(363,34){7}
//: {8}(98,139)(50,139){9}
reg c;    //: /sn:0 {0}(367,287)(104,287)(104,279){1}
//: {2}(106,277)(148,277){3}
//: {4}(102,277)(85,277){5}
//: {6}(83,275)(83,44)(363,44){7}
//: {8}(81,277)(52,277){9}
wire w6;    //: /sn:0 {0}(602,213)(602,229)(541,229){1}
wire w7;    //: /sn:0 {0}(157,356)(169,356){1}
//: {2}(173,356)(362,356){3}
//: {4}(171,354)(171,292)(367,292){5}
wire w16;    //: /sn:0 {0}(388,284)(406,284)(406,232)(520,232){1}
wire w19;    //: /sn:0 {0}(383,348)(420,348)(420,237)(520,237){1}
wire w3;    //: /sn:0 {0}(362,346)(205,346)(205,207)(174,207){1}
//: {2}(170,207)(160,207){3}
//: {4}(172,209)(172,282)(367,282){5}
wire w1;    //: /sn:0 {0}(362,341)(216,341)(216,141){1}
//: {2}(218,139)(242,139)(242,172)(368,172){3}
//: {4}(214,139)(158,139){5}
wire w8;    //: /sn:0 {0}(384,41)(485,41)(485,222)(520,222){1}
wire w13;    //: /sn:0 {0}(389,179)(423,179)(423,227)(520,227){1}
wire w5;    //: /sn:0 {0}(368,182)(240,182)(240,277)(183,277){1}
//: {2}(179,277)(164,277){3}
//: {4}(181,279)(181,351)(362,351){5}
//: enddecls

  //: joint g8 (a) @(112, 139) /w:[ 4 6 3 -1 ]
  _GGNBUF #(2) g4 (.I(a), .Z(w1));   //: @(148,139) /sn:0 /w:[ 5 5 ]
  _GGAND4 #(10) g13 (.I0(a), .I1(w3), .I2(c), .I3(w7), .Z(w16));   //: @(378,284) /sn:0 /w:[ 0 5 0 5 0 ]
  //: SWITCH g3 (d) @(32,356) /sn:0 /w:[ 9 ] /st:0 /dn:1
  //: SWITCH g2 (c) @(35,277) /sn:0 /w:[ 9 ] /st:0 /dn:1
  //: SWITCH g1 (b) @(30,207) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g16 (c) @(83, 277) /w:[ 5 6 8 -1 ]
  _GGAND4 #(10) g11 (.I0(a), .I1(b), .I2(c), .I3(d), .Z(w8));   //: @(374,41) /sn:0 /w:[ 7 9 7 3 0 ]
  _GGOR4 #(10) g10 (.I0(w8), .I1(w13), .I2(w16), .I3(w19), .Z(w6));   //: @(531,229) /sn:0 /w:[ 1 1 1 1 1 ]
  //: joint g19 (w5) @(181, 277) /w:[ 1 -1 2 4 ]
  _GGNBUF #(2) g6 (.I(c), .Z(w5));   //: @(154,277) /sn:0 /w:[ 3 3 ]
  //: LED g9 (w6) @(602,206) /sn:0 /w:[ 0 ] /type:0
  _GGNBUF #(2) g7 (.I(d), .Z(w7));   //: @(147,356) /sn:0 /w:[ 7 0 ]
  //: joint g20 (b) @(91, 178) /w:[ 6 8 -1 5 ]
  //: joint g15 (b) @(91, 207) /w:[ 2 4 1 -1 ]
  //: joint g25 (c) @(104, 277) /w:[ 2 -1 4 1 ]
  //: joint g17 (d) @(72, 356) /w:[ 6 5 8 -1 ]
  _GGAND4 #(10) g14 (.I0(w1), .I1(w3), .I2(w5), .I3(w7), .Z(w19));   //: @(373,348) /sn:0 /w:[ 0 0 5 3 0 ]
  _GGNBUF #(2) g5 (.I(b), .Z(w3));   //: @(150,207) /sn:0 /w:[ 3 3 ]
  //: joint g24 (a) @(100, 139) /w:[ 2 -1 8 1 ]
  //: joint g21 (d) @(72, 187) /w:[ 1 2 -1 4 ]
  //: joint g23 (w3) @(172, 207) /w:[ 1 -1 2 4 ]
  //: joint g22 (w7) @(171, 356) /w:[ 2 4 1 -1 ]
  //: SWITCH g0 (a) @(33,139) /sn:0 /w:[ 9 ] /st:0 /dn:1
  //: joint g18 (w1) @(216, 139) /w:[ 2 -1 4 1 ]
  _GGAND4 #(10) g12 (.I0(w1), .I1(b), .I2(w5), .I3(d), .Z(w13));   //: @(379,179) /sn:0 /w:[ 3 7 0 0 0 ]

endmodule
//: /netlistEnd

